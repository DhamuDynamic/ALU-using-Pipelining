// ALU Design using Pipelining
module ALU(clk1,clk2,rs1,rs2,rd,addr,func,y);
	input clk1,clk2;
	input [3:0] rs1,rs2,rd,func;
	input [7:0] addr;
	output [15:0] y;
	reg [15:0] L12_A,L12_B,L23_y,L34_y;
	reg [3:0] L12_rd,L12_func,L23_rd;
	reg [7:0] L12_addr,L23_addr,L34_addr;
	reg [15:0] RegBank [0:15];
	reg [15:0] Mem [0:255];
	assign y = L34_y;
	always @(posedge clk1)
		begin
			L12_A <= #2 RegBank[rs1];
			L12_B <= #2 RegBank[rs2];
			L12_rd <= #2 rd;
			L12_func <= #2 func;
			L12_addr <= addr;
		end
	always @(negedge clk2)
		begin
			case(func)
				0 : L23_y <= #2 L12_A + L12_B;
				1 : L23_y <= #2 L12_A - L12_B;
				2 : L23_y <= #2 L12_A * L12_B;
				3 : L23_y <= #2 L12_A;
				4 : L23_y <= #2 L12_B;
				5 : L23_y <= #2 L12_A & L12_B;
				6 : L23_y <= #2 L12_A | L12_B;
				7 : L23_y <= #2 L12_A ^ L12_B;
				8 : L23_y <= #2 L12_A >> 1;
				9 : L23_y <= #2 L12_A << 1;
				10 : L23_y <= #2 L12_B >> 1;
				default : L23_y <= #2 16'hx;
			endcase
			L23_rd <= #2 L12_rd;
			L23_addr <= L23_addr;
		end
	always @(posedge clk1)
		begin
			RegBank[L23_rd] <= #2 L23_y;
			L34_y <= #2 L23_y;
			L34_addr <= L23_addr;
		end
	always @(negedge clk2)
		begin
			Mem[L34_addr] <= #2 L34_y;
		end
endmodule
